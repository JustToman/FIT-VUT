-- fsm.vhd: Finite State Machine
-- Author(s): 
--
library ieee;
use ieee.std_logic_1164.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity fsm is
port(
   CLK         : in  std_logic;
   RESET       : in  std_logic;

   -- Input signals
   KEY         : in  std_logic_vector(15 downto 0);
   CNT_OF      : in  std_logic;

   -- Output signals
   FSM_CNT_CE  : out std_logic;
   FSM_MX_MEM  : out std_logic;
   FSM_MX_LCD  : out std_logic;
   FSM_LCD_WR  : out std_logic;
   FSM_LCD_CLR : out std_logic
);
end entity fsm;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture behavioral of fsm is
   type t_state is (TEST1,TEST2,TEST3,TEST4,TEST5,TEST16,TEST17,TEST18,TEST19,TEST110,TEST111,TEST26,TEST27,TEST28,TEST29,TEST210,TEST_ERR,TEST_OK,PRINT_OK,PRINT_ERROR, FINISH);
   signal present_state, next_state : t_state;

begin 
-- -------------------------------------------------------
sync_logic : process(RESET, CLK)
begin
   if (RESET = '1') then
      present_state <= TEST1;
   elsif (CLK'event AND CLK = '1') then
      present_state <= next_state;
   end if;
end process sync_logic;

-- -------------------------------------------------------
next_state_logic : process(present_state, KEY, CNT_OF)
begin
   case (present_state) is
	-- - - - - - - - - - - - - - - - - - - - - - -
   when TEST1 =>
		next_state <= TEST1;
      if (KEY(1) = '1') then 
			next_state <= TEST2;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR; 
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
   when TEST2 =>
		next_state <= TEST2;
      if (KEY(4) = '1') then 
			next_state <= TEST3;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR; 
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST3 =>
		next_state <= TEST3;
      if (KEY(9) = '1') then 
			next_state <= TEST4;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;   
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST4 =>
		next_state <= TEST4;
      if (KEY(1) = '1') then 
			next_state <= TEST5;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR; 
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST5 =>
		next_state <= TEST5;
      if (KEY(7) = '1') then 
			next_state <= TEST16;
		elsif (KEY(6) = '1') then 
			next_state <= TEST26; 
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST16 =>
		next_state <= TEST16;
      if (KEY(8) = '1') then 
			next_state <= TEST17;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST17 =>
		next_state <= TEST17;
      if (KEY(5) = '1') then 
			next_state <= TEST18;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR; 
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST18 =>
		next_state <= TEST18;
      if (KEY(8) = '1') then 
			next_state <= TEST19;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR; 
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST19 =>
		next_state <= TEST19;
      if (KEY(8) = '1') then 
			next_state <= TEST110;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR; 
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST110 =>
		next_state <= TEST110;
      if (KEY(1) = '1') then 
			next_state <= TEST111;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST111 =>
		next_state <= TEST111;
      if (KEY(6) = '1') then 
			next_state <= TEST_OK;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST26 =>
		next_state <= TEST26 ;
      if (KEY(1) = '1') then 
			next_state <= TEST27;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST27 =>
		next_state <= TEST27;
      if (KEY(9) = '1') then 
			next_state <= TEST28;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST28 =>
		next_state <= TEST28;
      if (KEY(6) = '1') then 
			next_state <= TEST29;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST29 =>
		next_state <= TEST29;
      if (KEY(0) = '1') then 
			next_state <= TEST210;
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST210 =>
		next_state <= TEST210;
      if (KEY(5) = '1') then 
			next_state <= TEST_OK; 
		elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_ERROR;  
      end if;
	-- - - - - - - - - - - - - - - - - - - - - - -
	 when TEST_ERR =>
		next_state <= TEST_ERR;
      if (KEY(15) = '1') then
         next_state <= PRINT_ERROR;
      end if;
	-- - ----- - - - - - - - - - - - - - - - - - - 
	when TEST_OK =>
		next_state <= TEST_OK;
      if (KEY(14 downto 0) /= "000000000000000") then
			next_state <= TEST_ERR;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_OK;
      end if;

   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_OK =>
      next_state <= PRINT_OK;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_ERROR =>
      next_state <= PRINT_ERROR;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when FINISH =>
      next_state <= FINISH;
      if (KEY(15) = '1') then
         next_state <= TEST1; 
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
      next_state <= TEST1;
   end case;
end process next_state_logic;

-- -------------------------------------------------------
output_logic : process(present_state, KEY)
begin
   FSM_CNT_CE     <= '0';
   FSM_MX_MEM     <= '0';
   FSM_MX_LCD     <= '0';
   FSM_LCD_WR     <= '0';
   FSM_LCD_CLR    <= '0';

   case (present_state) is
   -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST1 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST2 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST3 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST4 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST5 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST16 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST17 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST18 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST19 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST110 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	 -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST111 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	when TEST26 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	when TEST27 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	when TEST28 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	when TEST29 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	when TEST210 =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	when TEST_ERR | TEST_OK =>
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
	
   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_ERROR =>
		FSM_MX_MEM     <= '0';
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_LCD_WR     <= '1';
	 
	 when PRINT_OK =>
		FSM_MX_MEM     <= '1';
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_LCD_WR     <= '1';
      
   when FINISH =>
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
   end case;
end process output_logic;

end architecture behavioral;

